
`include "interface.sv"
`include "common.sv"
`include "transaction.sv"
`include "bfm.sv"
`include "generator.sv"
`include "agent.sv"
`include "env.sv"
`include "program.sv"
