program count_pro();
  
  count_env env;
  
  initial begin
    env=new();
    env.run();
  end
  
endprogram