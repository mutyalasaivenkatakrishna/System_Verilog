`include "memory.v"
`include "interface.sv"
`include "common.sv"
`include "mem_assert.sv"
`include "tx.sv"
`include "bfm.sv"
`include "gen.sv"
`include "monitor.sv"
`include "coverage.sv"
`include "score_board.sv"
`include "agent.sv"
`include "env.sv"
`include "top.sv"


// Open the files in the Order as follows for the better Understanding

// top.sv

//// agent.sv   ( jst see once )
//// env.sv     ( jst see once )

// interface.sv
// common.sv
// tx.sv
// gen.sv
// bfm.sv

// monitor.sv

// score_board.sv

// coverage.sv

// mem_assert.sv
// agent.sv
// env.sv
